dff d flip flop parametrized width default of 1 module dff d clk q parameter width 1 input clk input width 1 0 d output width 1 0 q reg width 1 0 q always posedge clk q d endmodule dffr d flip flop with active high synchronous reset parametrized width default of 1 module dffr d r clk q parameter width 1 input r input clk input width 1 0 d output width 1 0 q reg width 1 0 q always posedge clk if r q width 1 b0 else q d endmodule dffre d flip flop with active high enable and reset parametrized width default of 1 module dffre d en r clk q parameter width 1 input en input r input clk input width 1 0 d output width 1 0 q reg width 1 0 q always posedge clk if r q width 1 b0 else if en q d else q q endmodule
